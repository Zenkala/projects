library ieee;
use ieee.std_logic_1164.all;

entity pwm_gen is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity pwm_gen;

architecture RTL of pwm_gen is
	
begin

end architecture RTL;
